module microprocessorController();
endmodule
